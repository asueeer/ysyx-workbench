module shifter(
	input clk,
	output reg [7:0] Q);
	

endmodule
